module router #(
	parameter
)(

);
	

endmodule
