module dmux24(
    input [1:0]         s,
    output reg [3:0]    y
);
    always @(*) begin
        case(s)
            2'd0: y = 4'b0001;
            2'd1: y = 4'b0010;
            2'd2: y = 4'b0100;
            2'd2: y = 4'b1000;
        endcase
    end
endmodule