module sum (input x, y, output z);
    assign z = x + y;
endmodule // sum (input x, output y)